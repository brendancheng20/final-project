module bitwise_and(in1, in2, result);

	input[31:0] in1, in2;
	output[31:0] result;
	
	and and0(result[0], in1[0], in2[0]);
	and and1(result[1], in1[1], in2[1]);
	and and2(result[2], in1[2], in2[2]);
	and and3(result[3], in1[3], in2[3]);
	and and4(result[4], in1[4], in2[4]);
	and and5(result[5], in1[5], in2[5]);
	and and6(result[6], in1[6], in2[6]);
	and and7(result[7], in1[7], in2[7]);
	and and8(result[8], in1[8], in2[8]);
	and and9(result[9], in1[9], in2[9]);
	and and10(result[10], in1[10], in2[10]);
	and and11(result[11], in1[11], in2[11]);
	and and12(result[12], in1[12], in2[12]);
	and and13(result[13], in1[13], in2[13]);
	and and14(result[14], in1[14], in2[14]);
	and and15(result[15], in1[15], in2[15]);
	and and16(result[16], in1[16], in2[16]);
	and and17(result[17], in1[17], in2[17]);
	and and18(result[18], in1[18], in2[18]);
	and and19(result[19], in1[19], in2[19]);
	and and20(result[20], in1[20], in2[20]);
	and and21(result[21], in1[21], in2[21]);
	and and22(result[22], in1[22], in2[22]);
	and and23(result[23], in1[23], in2[23]);
	and and24(result[24], in1[24], in2[24]);
	and and25(result[25], in1[25], in2[25]);
	and and26(result[26], in1[26], in2[26]);
	and and27(result[27], in1[27], in2[27]);
	and and28(result[28], in1[28], in2[28]);
	and and29(result[29], in1[29], in2[29]);
	and and30(result[30], in1[30], in2[30]);
	and and31(result[31], in1[31], in2[31]);
	
endmodule
